library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;
use work.all;
use work.bus_multiplexer_pkg.all;

-- Testbench Processor Adiabatic Bifurcation

entity tb is
end entity tb;

architecture test of tb is

	component NSpinSolver is
		generic	(
				INT 					: integer := 5;
				FRAC					: integer := 9;
				M						: integer := 2; -- Address lenght
				NSPIN					: integer := 3; -- Number of Spin
				N						: integer := 20; --Bits for iteration
				N_ITERATION				: integer := 1000 -- Number of iteration
				);
		port	(
				clk						: in std_logic;
				reset					: in std_logic;
				start					: in std_logic;
				Data_in					: in std_logic_vector(INT+FRAC-1 downto 0);
				done					: out std_logic;
				xReady					: out std_logic;
				yReady					: out std_logic;
				S						: out std_logic_vector(NSPIN-1 downto 0);
				X_out					: out bus_array(NSPIN-1 downto 0, INT+FRAC-1 downto 0);	
				Y_out					: out bus_array(NSPIN-1 downto 0, INT+FRAC-1 downto 0)
				);
	end component NSpinSolver;
	
	component clock_gen 
		port ( 
			  clk   : out std_logic
			  );
	end component clock_gen;
	
	
	file ParamFile, file_outputS, file_output_X_Y	: text;
	file ParamFileRandom							: text;
	signal clk										: std_logic;
	signal reset									: std_logic;
	signal start									: std_logic;
	signal done										: std_logic;
	signal xReady									: std_logic;
	signal yReady									: std_logic;
	
	signal data_in									: std_logic_vector(31 downto 0);
	signal X_out									: bus_array(49 downto 0, 31 downto 0);
	signal Y_out									: bus_array(49 downto 0, 31 downto 0);
	signal S										: std_logic_vector(49 downto 0);
	signal X0										: std_logic_vector(31 downto 0);
	signal Y0										: std_logic_vector(31 downto 0);
	signal S0										: std_logic;
	signal X1										: std_logic_vector(31 downto 0);
	signal Y1										: std_logic_vector(31 downto 0);
	signal S1										: std_logic;
	signal X2										: std_logic_vector(31 downto 0);
	signal Y2										: std_logic_vector(31 downto 0);
	signal S2										: std_logic;
	signal X3										: std_logic_vector(31 downto 0);
	signal Y3										: std_logic_vector(31 downto 0);
	signal S3										: std_logic;
	signal X4										: std_logic_vector(31 downto 0);
	signal Y4										: std_logic_vector(31 downto 0);
	signal S4										: std_logic;
	signal X5										: std_logic_vector(31 downto 0);
	signal Y5										: std_logic_vector(31 downto 0);
	signal S5										: std_logic;
	signal X6										: std_logic_vector(31 downto 0);
	signal Y6										: std_logic_vector(31 downto 0);
	signal S6										: std_logic;
	signal X7										: std_logic_vector(31 downto 0);
	signal Y7										: std_logic_vector(31 downto 0);
	signal S7										: std_logic;
	signal X8										: std_logic_vector(31 downto 0);
	signal Y8										: std_logic_vector(31 downto 0);
	signal S8										: std_logic;
	signal X9										: std_logic_vector(31 downto 0);
	signal Y9										: std_logic_vector(31 downto 0);
	signal S9										: std_logic;
	signal X10										: std_logic_vector(31 downto 0);
	signal Y10										: std_logic_vector(31 downto 0);
	signal S10										: std_logic;
	signal X11										: std_logic_vector(31 downto 0);
	signal Y11										: std_logic_vector(31 downto 0);
	signal S11										: std_logic;
	signal X12										: std_logic_vector(31 downto 0);
	signal Y12										: std_logic_vector(31 downto 0);
	signal S12										: std_logic;
	signal X13										: std_logic_vector(31 downto 0);
	signal Y13										: std_logic_vector(31 downto 0);
	signal S13										: std_logic;
	signal X14										: std_logic_vector(31 downto 0);
	signal Y14										: std_logic_vector(31 downto 0);
	signal S14										: std_logic;
	signal X15										: std_logic_vector(31 downto 0);
	signal Y15										: std_logic_vector(31 downto 0);
	signal S15										: std_logic;
	signal X16										: std_logic_vector(31 downto 0);
	signal Y16										: std_logic_vector(31 downto 0);
	signal S16										: std_logic;
	signal X17										: std_logic_vector(31 downto 0);
	signal Y17										: std_logic_vector(31 downto 0);
	signal S17										: std_logic;
	signal X18										: std_logic_vector(31 downto 0);
	signal Y18										: std_logic_vector(31 downto 0);
	signal S18										: std_logic;
	signal X19										: std_logic_vector(31 downto 0);
	signal Y19										: std_logic_vector(31 downto 0);
	signal S19										: std_logic;
	signal X20										: std_logic_vector(31 downto 0);
	signal Y20										: std_logic_vector(31 downto 0);
	signal S20										: std_logic;
	signal X21										: std_logic_vector(31 downto 0);
	signal Y21										: std_logic_vector(31 downto 0);
	signal S21										: std_logic;
	signal X22										: std_logic_vector(31 downto 0);
	signal Y22										: std_logic_vector(31 downto 0);
	signal S22										: std_logic;
	signal X23										: std_logic_vector(31 downto 0);
	signal Y23										: std_logic_vector(31 downto 0);
	signal S23										: std_logic;
	signal X24										: std_logic_vector(31 downto 0);
	signal Y24										: std_logic_vector(31 downto 0);
	signal S24										: std_logic;
	signal X25										: std_logic_vector(31 downto 0);
	signal Y25										: std_logic_vector(31 downto 0);
	signal S25										: std_logic;
	signal X26										: std_logic_vector(31 downto 0);
	signal Y26										: std_logic_vector(31 downto 0);
	signal S26										: std_logic;
	signal X27										: std_logic_vector(31 downto 0);
	signal Y27										: std_logic_vector(31 downto 0);
	signal S27										: std_logic;
	signal X28										: std_logic_vector(31 downto 0);
	signal Y28										: std_logic_vector(31 downto 0);
	signal S28										: std_logic;
	signal X29										: std_logic_vector(31 downto 0);
	signal Y29										: std_logic_vector(31 downto 0);
	signal S29										: std_logic;
	signal X30										: std_logic_vector(31 downto 0);
	signal Y30										: std_logic_vector(31 downto 0);
	signal S30										: std_logic;
	signal X31										: std_logic_vector(31 downto 0);
	signal Y31										: std_logic_vector(31 downto 0);
	signal S31										: std_logic;
	signal X32										: std_logic_vector(31 downto 0);
	signal Y32										: std_logic_vector(31 downto 0);
	signal S32										: std_logic;
	signal X33										: std_logic_vector(31 downto 0);
	signal Y33										: std_logic_vector(31 downto 0);
	signal S33										: std_logic;
	signal X34										: std_logic_vector(31 downto 0);
	signal Y34										: std_logic_vector(31 downto 0);
	signal S34										: std_logic;
	signal X35										: std_logic_vector(31 downto 0);
	signal Y35										: std_logic_vector(31 downto 0);
	signal S35										: std_logic;
	signal X36										: std_logic_vector(31 downto 0);
	signal Y36										: std_logic_vector(31 downto 0);
	signal S36										: std_logic;
	signal X37										: std_logic_vector(31 downto 0);
	signal Y37										: std_logic_vector(31 downto 0);
	signal S37										: std_logic;
	signal X38										: std_logic_vector(31 downto 0);
	signal Y38										: std_logic_vector(31 downto 0);
	signal S38										: std_logic;
	signal X39										: std_logic_vector(31 downto 0);
	signal Y39										: std_logic_vector(31 downto 0);
	signal S39										: std_logic;
	signal X40										: std_logic_vector(31 downto 0);
	signal Y40										: std_logic_vector(31 downto 0);
	signal S40										: std_logic;
	signal X41										: std_logic_vector(31 downto 0);
	signal Y41										: std_logic_vector(31 downto 0);
	signal S41										: std_logic;
	signal X42										: std_logic_vector(31 downto 0);
	signal Y42										: std_logic_vector(31 downto 0);
	signal S42										: std_logic;
	signal X43										: std_logic_vector(31 downto 0);
	signal Y43										: std_logic_vector(31 downto 0);
	signal S43										: std_logic;
	signal X44										: std_logic_vector(31 downto 0);
	signal Y44										: std_logic_vector(31 downto 0);
	signal S44										: std_logic;
	signal X45										: std_logic_vector(31 downto 0);
	signal Y45										: std_logic_vector(31 downto 0);
	signal S45										: std_logic;
	signal X46										: std_logic_vector(31 downto 0);
	signal Y46										: std_logic_vector(31 downto 0);
	signal S46										: std_logic;
	signal X47										: std_logic_vector(31 downto 0);
	signal Y47										: std_logic_vector(31 downto 0);
	signal S47										: std_logic;
	signal X48										: std_logic_vector(31 downto 0);
	signal Y48										: std_logic_vector(31 downto 0);
	signal S48										: std_logic;
	signal X49										: std_logic_vector(31 downto 0);
	signal Y49										: std_logic_vector(31 downto 0);
	signal S49										: std_logic;

	
	begin
	
		DUT : NSpinSolver
					generic map (
		
								INT 					=> 12,
								FRAC 					=> 20,
								M 					    => 6,
								NSPIN 					=> 50,
								N 					    => 8,
								N_ITERATION	 		=> 200
								)
					port map	(
								clk						=> clk,
								reset					=> reset,
								start					=> start,
								Data_in					=> data_in,
								done					=> done, 
								xReady					=> xReady,
								yReady					=> yReady,
								S						=> S, 
								X_out					=> X_out,
								Y_out					=> Y_out
								);
		slv_from_slm_row(X0, X_out, 0);
		slv_from_slm_row(Y0, Y_out, 0);
		S0					<= S(0);
		slv_from_slm_row(X1, X_out, 1);
		slv_from_slm_row(Y1, Y_out, 1);
		S1					<= S(1);
		slv_from_slm_row(X2, X_out, 2);
		slv_from_slm_row(Y2, Y_out, 2);
		S2					<= S(2);
		slv_from_slm_row(X3, X_out, 3);
		slv_from_slm_row(Y3, Y_out, 3);
		S3					<= S(3);
		slv_from_slm_row(X4, X_out, 4);
		slv_from_slm_row(Y4, Y_out, 4);
		S4					<= S(4);
		slv_from_slm_row(X5, X_out, 5);
		slv_from_slm_row(Y5, Y_out, 5);
		S5					<= S(5);
		slv_from_slm_row(X6, X_out, 6);
		slv_from_slm_row(Y6, Y_out, 6);
		S6					<= S(6);
		slv_from_slm_row(X7, X_out, 7);
		slv_from_slm_row(Y7, Y_out, 7);
		S7					<= S(7);
		slv_from_slm_row(X8, X_out, 8);
		slv_from_slm_row(Y8, Y_out, 8);
		S8					<= S(8);
		slv_from_slm_row(X9, X_out, 9);
		slv_from_slm_row(Y9, Y_out, 9);
		S9					<= S(9);
		slv_from_slm_row(X10, X_out, 10);
		slv_from_slm_row(Y10, Y_out, 10);
		S10					<= S(10);
		slv_from_slm_row(X11, X_out, 11);
		slv_from_slm_row(Y11, Y_out, 11);
		S11					<= S(11);
		slv_from_slm_row(X12, X_out, 12);
		slv_from_slm_row(Y12, Y_out, 12);
		S12					<= S(12);
		slv_from_slm_row(X13, X_out, 13);
		slv_from_slm_row(Y13, Y_out, 13);
		S13					<= S(13);
		slv_from_slm_row(X14, X_out, 14);
		slv_from_slm_row(Y14, Y_out, 14);
		S14					<= S(14);
		slv_from_slm_row(X15, X_out, 15);
		slv_from_slm_row(Y15, Y_out, 15);
		S15					<= S(15);
		slv_from_slm_row(X16, X_out, 16);
		slv_from_slm_row(Y16, Y_out, 16);
		S16					<= S(16);
		slv_from_slm_row(X17, X_out, 17);
		slv_from_slm_row(Y17, Y_out, 17);
		S17					<= S(17);
		slv_from_slm_row(X18, X_out, 18);
		slv_from_slm_row(Y18, Y_out, 18);
		S18					<= S(18);
		slv_from_slm_row(X19, X_out, 19);
		slv_from_slm_row(Y19, Y_out, 19);
		S19					<= S(19);
		slv_from_slm_row(X20, X_out, 20);
		slv_from_slm_row(Y20, Y_out, 20);
		S20					<= S(20);
		slv_from_slm_row(X21, X_out, 21);
		slv_from_slm_row(Y21, Y_out, 21);
		S21					<= S(21);
		slv_from_slm_row(X22, X_out, 22);
		slv_from_slm_row(Y22, Y_out, 22);
		S22					<= S(22);
		slv_from_slm_row(X23, X_out, 23);
		slv_from_slm_row(Y23, Y_out, 23);
		S23					<= S(23);
		slv_from_slm_row(X24, X_out, 24);
		slv_from_slm_row(Y24, Y_out, 24);
		S24					<= S(24);
		slv_from_slm_row(X25, X_out, 25);
		slv_from_slm_row(Y25, Y_out, 25);
		S25					<= S(25);
		slv_from_slm_row(X26, X_out, 26);
		slv_from_slm_row(Y26, Y_out, 26);
		S26					<= S(26);
		slv_from_slm_row(X27, X_out, 27);
		slv_from_slm_row(Y27, Y_out, 27);
		S27					<= S(27);
		slv_from_slm_row(X28, X_out, 28);
		slv_from_slm_row(Y28, Y_out, 28);
		S28					<= S(28);
		slv_from_slm_row(X29, X_out, 29);
		slv_from_slm_row(Y29, Y_out, 29);
		S29					<= S(29);
		slv_from_slm_row(X30, X_out, 30);
		slv_from_slm_row(Y30, Y_out, 30);
		S30					<= S(30);
		slv_from_slm_row(X31, X_out, 31);
		slv_from_slm_row(Y31, Y_out, 31);
		S31					<= S(31);
		slv_from_slm_row(X32, X_out, 32);
		slv_from_slm_row(Y32, Y_out, 32);
		S32					<= S(32);
		slv_from_slm_row(X33, X_out, 33);
		slv_from_slm_row(Y33, Y_out, 33);
		S33					<= S(33);
		slv_from_slm_row(X34, X_out, 34);
		slv_from_slm_row(Y34, Y_out, 34);
		S34					<= S(34);
		slv_from_slm_row(X35, X_out, 35);
		slv_from_slm_row(Y35, Y_out, 35);
		S35					<= S(35);
		slv_from_slm_row(X36, X_out, 36);
		slv_from_slm_row(Y36, Y_out, 36);
		S36					<= S(36);
		slv_from_slm_row(X37, X_out, 37);
		slv_from_slm_row(Y37, Y_out, 37);
		S37					<= S(37);
		slv_from_slm_row(X38, X_out, 38);
		slv_from_slm_row(Y38, Y_out, 38);
		S38					<= S(38);
		slv_from_slm_row(X39, X_out, 39);
		slv_from_slm_row(Y39, Y_out, 39);
		S39					<= S(39);
		slv_from_slm_row(X40, X_out, 40);
		slv_from_slm_row(Y40, Y_out, 40);
		S40					<= S(40);
		slv_from_slm_row(X41, X_out, 41);
		slv_from_slm_row(Y41, Y_out, 41);
		S41					<= S(41);
		slv_from_slm_row(X42, X_out, 42);
		slv_from_slm_row(Y42, Y_out, 42);
		S42					<= S(42);
		slv_from_slm_row(X43, X_out, 43);
		slv_from_slm_row(Y43, Y_out, 43);
		S43					<= S(43);
		slv_from_slm_row(X44, X_out, 44);
		slv_from_slm_row(Y44, Y_out, 44);
		S44					<= S(44);
		slv_from_slm_row(X45, X_out, 45);
		slv_from_slm_row(Y45, Y_out, 45);
		S45					<= S(45);
		slv_from_slm_row(X46, X_out, 46);
		slv_from_slm_row(Y46, Y_out, 46);
		S46					<= S(46);
		slv_from_slm_row(X47, X_out, 47);
		slv_from_slm_row(Y47, Y_out, 47);
		S47					<= S(47);
		slv_from_slm_row(X48, X_out, 48);
		slv_from_slm_row(Y48, Y_out, 48);
		S48					<= S(48);
		slv_from_slm_row(X49, X_out, 49);
		slv_from_slm_row(Y49, Y_out, 49);
		S49					<= S(49);
								
		clkGen: clock_gen 
					port  map	( 
								clk					=> clk
								);
								
							
		read_files_process: process
									variable v_ILINEP    		: line;
									variable v_ILINEYR    		: line;
									variable v_OLINE    		: line;
									variable v_OLINE_X_Y    	: line;
									variable i 					: integer := 0;
									variable k 					: integer := 0;
									variable y 					: integer := 0;
									variable space 				: character;
			
									variable data_in_v 			: std_logic_vector(31 downto 0);
									begin
									file_open(ParamFileRandom, "resultsMaxCut1/Problem_50_y_init_variables.txt", read_mode);
									file_open(file_outputS, "resultsMaxCut1/output_file_50.txt", write_mode);
									file_open(file_output_X_Y, "resultsMaxCut1/output_file_X_Y_50.txt", write_mode);
									while i < 1 loop
										start <= '0';
										reset <= '0';
										wait for 12 ns;
										reset <= '1';
										wait for 12 ns;
										start <= '1';
										wait for 10 ns;
										start <= '0';
										k := 0;
								
										file_open(ParamFile, "resultsMaxCut1/InputParameter_50.txt", read_mode);
								
									while not endfile(ParamFile) loop
										-- read the parameters
										-- We read in order the following parameters:
										-- ShapePt, Delta4K, K_1, offset, Delta, xi
										-- deltaT, HVector0, HVector1, J12, J21, YOld
										if k = 56 then
											readline(ParamFileRandom, v_ILINEYR);
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											read(v_ILINEYR, space);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
											read(v_ILINEYR, y);
											data_in <= std_logic_vector(to_signed(y, 32));
											wait for 10 ns;
										else
											readline(ParamFile, v_ILINEP);
											read(v_ILINEP, data_in_v);
											data_in <= data_in_v;
											wait for 10 ns;
										end if;
										k:= k+1;
										
									end loop;
									--close parameters file
									file_close(ParamFile);
									loop
										wait until xReady = '1' or done ='1';
										if done = '1' then
											exit;
										end if;
										wait for 12 ns;
										write(v_OLINE_X_Y, X0);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X1);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X2);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X3);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X4);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X5);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X6);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X7);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X8);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X9);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X10);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X11);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X12);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X13);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X14);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X15);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X16);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X17);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X18);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X19);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X20);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X21);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X22);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X23);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X24);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X25);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X26);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X27);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X28);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X29);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X30);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X31);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X32);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X33);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X34);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X35);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X36);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X37);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X38);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X39);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X40);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X41);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X42);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X43);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X44);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X45);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X46);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X47);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X48);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, X49);
										write(v_OLINE_X_Y, ' ');
										wait until yReady = '1';
										wait for 8 ns;
										write(v_OLINE_X_Y, Y0);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y1);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y2);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y3);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y4);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y5);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y6);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y7);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y8);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y9);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y10);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y11);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y12);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y13);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y14);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y15);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y16);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y17);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y18);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y19);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y20);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y21);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y22);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y23);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y24);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y25);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y26);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y27);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y28);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y29);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y30);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y31);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y32);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y33);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y34);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y35);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y36);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y37);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y38);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y39);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y40);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y41);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y42);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y43);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y44);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y45);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y46);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y47);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y48);
										write(v_OLINE_X_Y, ' ');
										write(v_OLINE_X_Y, Y49);
										writeline(file_output_X_Y, v_OLINE_X_Y);
									
									end loop;
					
	
									wait for 11 ns; -- wait for one clock period	
									write(v_OLINE, S0);
									write(v_OLINE, ' ');
									write(v_OLINE, S1);
									write(v_OLINE, ' ');
									write(v_OLINE, S2);
									write(v_OLINE, ' ');
									write(v_OLINE, S3);
									write(v_OLINE, ' ');
									write(v_OLINE, S4);
									write(v_OLINE, ' ');
									write(v_OLINE, S5);
									write(v_OLINE, ' ');
									write(v_OLINE, S6);
									write(v_OLINE, ' ');
									write(v_OLINE, S7);
									write(v_OLINE, ' ');
									write(v_OLINE, S8);
									write(v_OLINE, ' ');
									write(v_OLINE, S9);
									write(v_OLINE, ' ');
									write(v_OLINE, S10);
									write(v_OLINE, ' ');
									write(v_OLINE, S11);
									write(v_OLINE, ' ');
									write(v_OLINE, S12);
									write(v_OLINE, ' ');
									write(v_OLINE, S13);
									write(v_OLINE, ' ');
									write(v_OLINE, S14);
									write(v_OLINE, ' ');
									write(v_OLINE, S15);
									write(v_OLINE, ' ');
									write(v_OLINE, S16);
									write(v_OLINE, ' ');
									write(v_OLINE, S17);
									write(v_OLINE, ' ');
									write(v_OLINE, S18);
									write(v_OLINE, ' ');
									write(v_OLINE, S19);
									write(v_OLINE, ' ');
									write(v_OLINE, S20);
									write(v_OLINE, ' ');
									write(v_OLINE, S21);
									write(v_OLINE, ' ');
									write(v_OLINE, S22);
									write(v_OLINE, ' ');
									write(v_OLINE, S23);
									write(v_OLINE, ' ');
									write(v_OLINE, S24);
									write(v_OLINE, ' ');
									write(v_OLINE, S25);
									write(v_OLINE, ' ');
									write(v_OLINE, S26);
									write(v_OLINE, ' ');
									write(v_OLINE, S27);
									write(v_OLINE, ' ');
									write(v_OLINE, S28);
									write(v_OLINE, ' ');
									write(v_OLINE, S29);
									write(v_OLINE, ' ');
									write(v_OLINE, S30);
									write(v_OLINE, ' ');
									write(v_OLINE, S31);
									write(v_OLINE, ' ');
									write(v_OLINE, S32);
									write(v_OLINE, ' ');
									write(v_OLINE, S33);
									write(v_OLINE, ' ');
									write(v_OLINE, S34);
									write(v_OLINE, ' ');
									write(v_OLINE, S35);
									write(v_OLINE, ' ');
									write(v_OLINE, S36);
									write(v_OLINE, ' ');
									write(v_OLINE, S37);
									write(v_OLINE, ' ');
									write(v_OLINE, S38);
									write(v_OLINE, ' ');
									write(v_OLINE, S39);
									write(v_OLINE, ' ');
									write(v_OLINE, S40);
									write(v_OLINE, ' ');
									write(v_OLINE, S41);
									write(v_OLINE, ' ');
									write(v_OLINE, S42);
									write(v_OLINE, ' ');
									write(v_OLINE, S43);
									write(v_OLINE, ' ');
									write(v_OLINE, S44);
									write(v_OLINE, ' ');
									write(v_OLINE, S45);
									write(v_OLINE, ' ');
									write(v_OLINE, S46);
									write(v_OLINE, ' ');
									write(v_OLINE, S47);
									write(v_OLINE, ' ');
									write(v_OLINE, S48);
									write(v_OLINE, ' ');
									write(v_OLINE, S49);
									writeline(file_outputS, v_OLINE);
									write(v_OLINE_X_Y, '_');
									writeline(file_output_X_Y, v_OLINE_X_Y);
									i:=i+1;
									end loop;
									--close output file
									file_close(file_outputS);
									file_close(file_output_X_Y);	
									file_close(ParamFileRandom);
									wait;
							end process;
end architecture test;
